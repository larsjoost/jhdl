

module test (a, b);

endmodule // test

package ENV is
  procedure STOP (STATUS: INTEGER);
end package ENV;

package body ENV is

  procedure STOP (STATUS: INTEGER) is
  begin
  end;

end package body ENV;

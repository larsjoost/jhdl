
package test_pkg is

  constant c : integer := 2;

end package test_pkg;

use work.test_pkg.all;

entity test is
end entity test;

architecture rtl of test is
begin
end architecture rtl;

entity test is
end entfity test;

architecture rtl of test is
begin
end architecture rtl;

entity test is
end entity test;

architecture rtl of test is

  type test_t is range 1 to 20;

begin
end architecture rtl;

entity test is
end entfity test;



package test is

  constant c : integer := 10;
  
  function test_function (
    a : integer;
    b : integer)
    return integer;

end package test;

entity test is
end entity   badname;


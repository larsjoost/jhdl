
use lib.pack.all;

entity test is
end entity test;

architecture rtl of test is
begin
end architecture rtl;

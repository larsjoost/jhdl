

-- Test 2

entity test is
end entity test;

-- Test 3

architecture rtl of test is
begin
end architecture rtl;

entity test is
end entity test;

architecture rtl of test is

  type range_t is range 0 to 1.0;
  
begin

end architecture rtl;
